
/* ----------------------------------------------------------------------------------------------- //
Project Title: UVM-Based Functional Verification of PCIe PHY Layer
Institution: University of Science and Technology, Zewail City
Project Team: Marwan Eid - Alaa Taha - Pater Gad - Almomenbelah Allam - Mahmoud Marzouk
File Description: Tx ALU Package
Version: 1.0
// ----------------------------------------------------------------------------------------------- */

package ALU_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    
    `include "ALU_cfg_obj.svh"
    `include "ALU_sequence_item.svh"
    `include "ALU_sequence.svh"
    `include "ALU_sequencer.svh"
    `include "ALU_driver.svh"
    `include "ALU_monitor.svh"
    `include "ALU_agent.svh"
    `include "ALU_subscriber.svh"
    `include "ALU_scoreboard.svh"
    `include "ALU_env.svh"    
    `include "ALU_test_base_class.svh"
    `include "ALU_test.svh"
    
    
endpackage: ALU_pkg
