
`ifndef CYCLE 
  `define CYCLE 10 
`endif 
`ifndef Tdrive 
  `define Tdrive #(0.2*`CYCLE) 
`endif 
`timescale 1ns/1ps